`timescale 1ns / 1ps

module Shifter_2(
    input [31:0] Input,
    output [31:0] Output
    );
	 
	 assign Output = Input ;


endmodule
